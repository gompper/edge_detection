entity sobel is
	generic(
	
	);
	port(
		clk : in std_logic;
		reset: in std_logic;
	
	);
end entity sobel;